module Gray_to_Binary(OT,IN);
output [3:0]OT;
input [3:0]IN;

buf b1(OT[3],IN[3]);
xor xr1(OT[2],OT[3],IN[2]);
xor xr2(OT[1],OT[2],IN[1]);
xor xr3( OT[0],OT[1],IN[0]);

endmodule



module testgb;

reg [3:0]IN;
wire [3:0]OT;
Gray_to_Binary  g_b(OT,IN);

initial
begin

#0 IN = 4'd0;
#100 IN = 4'd1;
#100 IN = 4'd2;
#100 IN = 4'd3;
#100 IN = 4'd4;
end

endmodule                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
